entity top is
    i_sys_clk : in std_logic
end top;

architecture top_behav of top is
begin
    
end top_behav;